`timescale 1ns / 1ps

module NOT_Gate(input a, output y);
assign y=~(a);
endmodule

