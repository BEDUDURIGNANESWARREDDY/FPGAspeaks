`timescale 1ns / 1ps


module XOR_Gate(input a,b, output y);

assign y=a^b;
endmodule
